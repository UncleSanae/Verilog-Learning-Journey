module hello;
    initial begin
        $display("Hello World!My Verilog works XD");
        $finish;
    end
endmodule